`ifndef _defines_h_
`define _defines_h_

`define KEY_0 0
`define KEY_1 1
`define KEY_2 2
`define KEY_3 3
`define KEY_4 4
`define KEY_5 5
`define KEY_6 6
`define KEY_7 7
`define KEY_8 8
`define KEY_9 9
`define KEY_A 10
`define KEY_B 11
`define KEY_C 12
`define KEY_D 13
`define KEY_E 14
`define KEY_F 15
`define KEY_NONE 16

`define S_WPR 2'd0
`define S_OP  2'd1
`define S_OBL 2'd2
`define S_GON 2'd3

`define SL_A 3'd0
`define SL_B 3'd1

`define SL_ADD 3'd0
`define SL_SUB 3'd1
`define SL_XOR 3'd2
`define SL_OR  3'd3
`define SL_AND 3'd4

`define ASCII_A 8'h41
`define ASCII_B 8'h42
`define ASCII_D 8'h44
`define ASCII_N 8'h4e
`define ASCII_O 8'h4f
`define ASCII_R 8'h52
`define ASCII_S 8'h53
`define ASCII_U 8'h55
`define ASCII_X 8'h58

`endif